library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity hex_sedam_seg is
end hex_sedam_seg;

architecture Behavioral of hex_sedam_seg is

begin


end Behavioral;

